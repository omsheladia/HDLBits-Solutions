module top_module( output one );

// Insert your code here
    assign one = [fixme];

endmodule