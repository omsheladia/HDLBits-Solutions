module top_module( input in, output out );
    reg wr;
    assign wr = in;
    assign out = wr;

endmodule
